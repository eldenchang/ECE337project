// $Id: $
// File name:   tb_ff_add.sv
// Created:     12/1/2017
// Author:      Andrew Beatty
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: Testbench for Finite Field Addition Module.

module tb_ff_add ();

