// $Id: $
// File name:   tb_flexbyte_pts_sr.sv
// Created:     11/28/2017
// Author:      Andrew Beatty
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: Testbench for flexbyte_pts_sr.sv
